sample_id	BCL6_fusion	BCL2_fusion	MYC_fusion
